
LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.numeric_std.all;  



ENTITY DE10_TOP_LEVEL is
    PORT
    (
        MAX10_CLK1_50    :  IN  STD_LOGIC;
        KEY              :  IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
        SW               :  IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
        HEX0             :  OUT  STD_LOGIC_VECTOR(0 TO 6);
        HEX1             :  OUT  STD_LOGIC_VECTOR(0 TO 6);
        HEX2             :  OUT  STD_LOGIC_VECTOR(0 TO 6);
	GPIO_35           :  OUT STD_LOGIC;
	GPIO_34           :  IN STD_LOGIC;
	LEDR_8 : OUT STD_LOGIC
);
END entity DE10_TOP_LEVEL;

ARCHITECTURE RTL OF DE10_TOP_LEVEL IS 

    signal     rst, clk, trig, echo, led  : std_logic;
    signal distance_object : integer;
    signal    distance_unit, distance_dizaine, distance_centaine    :  integer;
    signal Echo_Pulse_Time : unsigned(21 downto 0);
    signal echo_pulse_state : std_logic;

BEGIN 
    echo <= GPIO_34;
    GPIO_35 <= trig;
    clk <= MAX10_CLK1_50;
    LEDR_8 <= led; 
   
TRIGGER : entity work.trigger port map(clk=>clk, trigger => trig);
MESURE_TEMPS_ECHO : entity work.MesureTempsEchoIN port map(echo_pulse=>echo, clk=>clk, Echo_Pulse_Time=>Echo_Pulse_Time, echo_pulse_state=>echo_pulse_state);
--MESURE_DISTANCE : entity work.MesureDistance port map(distance_object=>distance_object,echo_pulse_state=>echo_pulse_state,echo_pulse=>echo_pulse);
--CONVERT_DISTANCE : entity work.Convert_Distance port map(distance_centaine=>distance_centaine,distance_dizaine=>distance_dizaine,distance_unit=>distance_unit);


--ET5 : entity work.Convert_Distance_7seg port map(Distance_Unit => unities, Distance_Dizaine => tens, Distance_Centaine => hundreds);
SEVEN_SEG0 : entity work.Convert_Distance_7seg port map(Unit => HEX0);
SEVEN_SEG1 : entity work.Convert_Distance_7seg port map(Dizaine => HEX1);
SEVEN_SEG2 : entity work.Convert_Distance_7seg port map(Centaine => HEX2);



END architecture RTL;

